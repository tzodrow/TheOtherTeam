module spu();

endmodule