module sprite_mem_access(sprite_number, action, attribute_value, sprite_data, addr_a, addr_b, data_a, data_b);
	
endmodule