module ascii2hex(
		input [8:0] ascii,
		output [3:0] hex);
	
	case(ascii)
		
	endcase
	
endmodule