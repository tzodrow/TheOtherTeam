module instruction_fetch(
		input clk,
		input rst,
		input [21:0] pc,
		output [31:0] instr);
	
	
endmodule
		