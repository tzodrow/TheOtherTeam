module move_logic(input start, 
   input sprite_data_active, input sprite_data_moving, input[18:0] sprite_data_coord, input[7:0] sprite_data_image, input[7:0] sprite_data_speed,
   input[1:0] sprite_data_direction,    
   output draw_sprite_start, output sprite_data_re, output sprite_data_we, output[23:0] sprite_data_address, output[18:0] sprite_data_coord_write);







endmodule